module executor

// import os 

// TODO: implement semi auto mode logic