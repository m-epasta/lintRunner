module executor

